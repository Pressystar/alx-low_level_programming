b0VIM 8.1      �d�$.�  root                                    92fcfb7da80e                            ~root/alx-low_level_programming/0x15-file_io/100-elf_header.c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                     ��������m       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad  %   )     �       �  �  �  �  �  �  t  s  r  J     �  �  �  y  O    �  �  �  �  �  ~  _  >  :          �  �  �  �  �  y  w  C  9  7  5  3  /    �  �  �  �  �  �  �  |  {  O  M  L  ,  +      �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  p
  o
  T
  R
  ?
  -
  &
  
  
  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  s	  Q	  M	  %	  #	  	  	  �  �  �  �  �  �  �  �  s  K  D  ;  !      	    �  �  �  �  �  w  a  C  A  0        �  �  �  �  �  �  �  �  }  {  f  e  J  H  4      �  �  �  �  �  �  �  t  m  V  :  3       �  �  �  �  �  �  �  ~  b  [  R  8  $  "         �  �  �  �  �  �  �    c  B  -  )  (                                        */  * @e_type: Elf_type  * @e_ident: pointer to ELF type  * print_type - Entry point /** } e_ident[EI_ABIVERSION]); printf(" ABI Version: %d\n", { void print_abi(unsigned char *e_ident)  */  * @e_ident: The ELF Abi  * print_abi - Entry point /** } } e_ident[EI_OSABI]); printf("<unknown: %x>\n", default: break; printf("Standalone App\n"); case ELFOSABI_STANDALONE: break; printf("ARM\n"); case ELFOSABI_ARM: break; printf("UNIX - TRU64\n"); case ELFOSABI_TRU64: break; printf("UNIX - FreeBSD\n"); case ELFOSABI_FREEBSD: break; printf("UNIX - Solaris\n"); case ELFOSABI_SOLARIS: break; printf("UNIX - Linux\n"); case ELFOSABI_LINUX: break; printf("UNIX - NETBSD\n"); case ELFOSABI_NETBSD: break; printf("UNIX - HP-UX\n"); case ELFOSABI_HPUX: break; printf("UNIX - System V\n"); case ELFOSABI_NONE: { switch (e_ident[EI_OSABI])  printf(" OS/ABI: "); { void print_osabi(unsigned char *e_ident)  */  * @e_ident: pointer to ELF version  * print_osabi - Entry point /** } } break; printf("\n"); default: break; printf(" (current)\n"); case EV_CURRENT: { switch (e_ident[EI_VERSION]); e_ident[EI_VERSION]); printf(" Version: %d", { void print_version(unsigned char *e_ident)  */  * @e_ident: the pointer to ELF verson  * print_version - Entry point /** } } e_ident[EI_CLASS]); printf("<unknown: %x>\n", default: break; printf("2's complement, big endian\n"); case ELFDATA2MSB: break; printf("2's complement, little endian\n"); case ELFDATA2LSB: break; printf("none\n"); case ELFDATANONE: { switch(e_ident[EI_DATA])  printf(" Data: "); { void print_data(unsigned char *e_ident)  */  * @e_ident: pointer to ELF class  * print_data - Entry point /** } } e_ident([EI_CLASS])); printf("<unknown: %x>\n", default: break; printf("ELF64\n"); case ELFCLASS64: break; printf("ELF32\n"); case ELFCLASS32: break; printf("none\n"); case ELFCLASSNONE: { switch (e_ident[EI_CLASS])  printf(" Class: "); { void print_class(unsigned char *e_ident)  */  * @e_ident: ELF class  * print_class - Entry point /** } } printf(" "); else printf("\n"); if (index == EI_NIDENT - 1)  printf("%02x", e_ident[index]);  { for (index = 0; index < EI_NIDENT; index++)  printf(" Magic: ");  int index; { void print_magic(unsigned char *e_ident)  */  * Description: Magic numbers separated  * @e_ident: ELF magic numbers  * print_magic - Entry point /** } } } exit(98); dprintf(STDERR_FILENO, "Error: Not an ELF file\n"); { e_ident[index] != 'F') e_ident[index] != 'L' && e_ident[index] != 'E' && if (e_ident[index] != 127 && { for (index = 0; index < 4; index++)  int index; { void check_elf(unsigned char *e_ident)  */  * Description: negative exit 98  * @e_ident: elf magic numbers  * check_elf - write a function that checs file /**  void close_elf(int elf); unsigned char *e_ident); void print_entry(unsigned long int e_entry, void print_type(unsigned int e_type, unsigned char *e_ident); void print_osabi(unsigned char *e_ident); void print_abi(unsigned char *e_ident); void print_version(unsigned char *e_ident); void print_data(unsigned char *e_ident); void print_class(unsigned char *e_ident); void print_magic(unsigned char *e_ident); void check_elf(unsigned char *e_ident);   #include <stdlib.h> #include <stdio.h> #include <unistd.h> #include <fcntl.h> #include <sys/stat.h> #include <sys/types.h> #include <elf.h> ad  �  [     m       �  �  �  �  �  z  y  i  h  f  X  ?  8  +       �  �  �  �  �  �    a  Z  Q  .  ,  *  &  �  �  �  �  i  g  E  D      �  �  �  �  Z  U  :  8  4      �  �  �  �  �  �  n  d  b  `  \  F  (    �
  �
  �
  �
  �
  �
  v
  u
  X
  W
  J
  H
  	
  �	  �	  �	  �	  �	  �	  u	  k	  i	  @	  3	  1	  #	  	  �  �  �  �  �  w  Y  <    �  �  �  �  x  i  ]  [  Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             } return (0); close_elf(-o); free(header); print_entry(header->e_entry, header->e_ident); print_type(header->e_type, header->e_ident); print_abi(header->e_ident); print_osabi(header->e_ident); print_version(header->e_ident); print_data(header->e_ident); print_class(header->e_ident); print_magic(header->e_ident); printf("ELF Header:\n"); check_elf(header->e_ident); } exit(98); dprintf(STDERR_FILENO, "Error:'%s': No such file\n", argv[1]); close_elf(o); free(header); { if (r == -1) r = read(o, header, sizeof(Elf64_Ehdr)); } exit(98); dprintf(STDERR_FILENO, "Error:can't read file %s\n", argv[1]); close_elf(o); { if (header == NULL) header = malloc(sizeof(Elf64_Ehdr)); } exit(98); dprintf(STDERR_FILENO, "Error:Can't read file %s\n", argv[1]); { if (o == -1)  o = open(argv[1], O_RDONLY);  int o, r; Elf64_Ehdr *header; { int main(int __attribute__((__unused__))argc, char *argv[])  */  * Description:if negative exit code 98  * Return: 0  * @argv: array of arguments  * @argc: number of arguments  * main - Entry point /** } } exit(98); dprintf(STDERR_FILENO, "Error: Can't close fd %d\n", elf); { if (close(elf) == -1) { void close_elf(int elf)  */  * Description: can't close exit 98  * @elf: The ELF file  * close_elf - Entry point /** } printf("%#lx\n", e_entry); else printf("%#x\n", (unsigned int)e_entry); if (e_ident[EI_CLASS] == ELFCLASS32) } e_entry = (e_entry << 16) | (e_entry >> 16); e_entry = ((e_entry << 8) & 0xFF00FF00) | ((e_entry >> 8) & 0xFF00FF); { if (e_ident[EI_DATA] == ELFDATA2MSB)  printf(" Entry point address: "); { void print_entry(unsigned long int e_entry, unsigned char *e_ident)  */  * @e_ident: a pointer containing ELF class  * @e_entry: address  * print_entry - write a function that prints Entry /** } } printf("<unknown: %x>\n", e_type); default: break; printf("CORE (Core file)\n"); case ET_CORE: break; printf("DYN (Shared object file)\n"); case ET_DYN: break; printf("EXEC (Executable file)\n"); case ET_EXEC: break; printf("REL (Relocatable file)/n"); case ET_REL: break; printf("NONE (None)\n"); case ET_NONE: {  switch (e_type)  printf(" Type: ");  e_type >>= 8; if (e_ident[EI_DATA] == ELFDATA2MSB) { void print_type(unsigned int e_type, unsigned char *e_ident) 